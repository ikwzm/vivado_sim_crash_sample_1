-----------------------------------------------------------------------------------
--!     @file    aix4_test_1_2.vhd
--!     @brief   TEST BENCH No.1.2 for DUMMY_PLUG.AXI4_MODELS
--!     @version 1.5.0
--!     @date    2013/5/31
--!     @author  Ichiro Kawazome <ichiro_k@ca2.so-net.ne.jp>
-----------------------------------------------------------------------------------
--
--      Copyright (C) 2012,2013 Ichiro Kawazome
--      All rights reserved.
--
--      Redistribution and use in source and binary forms, with or without
--      modification, are permitted provided that the following conditions
--      are met:
--
--        1. Redistributions of source code must retain the above copyright
--           notice, this list of conditions and the following disclaimer.
--
--        2. Redistributions in binary form must reproduce the above copyright
--           notice, this list of conditions and the following disclaimer in
--           the documentation and/or other materials provided with the
--           distribution.
--
--      THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
--      "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
--      LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
--      A PARTICULAR PURPOSE ARE DISCLAIMED.  IN NO EVENT SHALL THE COPYRIGHT
--      OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
--      SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
--      LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
--      DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
--      THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT 
--      (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
--      OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--
-----------------------------------------------------------------------------------
library ieee;
use     ieee.std_logic_1164.all;
library DUMMY_PLUG;
use     DUMMY_PLUG.CORE.REPORT_STATUS_TYPE;
entity  DUMMY_PLUG_AXI4_TEST_1_2 is
end     DUMMY_PLUG_AXI4_TEST_1_2;
architecture MODEL of DUMMY_PLUG_AXI4_TEST_1_2 is
    constant NAME            : STRING  := "AXI4_TEST_1_2";
    constant SCENARIO_FILE   : STRING  := "../src/axi4_test_1_2.snr";
    constant EXP_REPORT      : REPORT_STATUS_TYPE := (
        valid          => TRUE,
        error_count    =>  0,
        mismatch_count =>  0,
        warning_count  =>  0,
        failure_count  =>  0
    );
    component DUMMY_PLUG_AXI4_TEST_1
        generic (
            NAME            : STRING;
            SCENARIO_FILE   : STRING;
            DATA_WIDTH      : integer;
            READ_ENABLE     : boolean;
            WRITE_ENABLE    : boolean;
            EXP_REPORT      : REPORT_STATUS_TYPE
        );
    end component;
begin
    U: DUMMY_PLUG_AXI4_TEST_1 generic map(NAME, SCENARIO_FILE, 64, TRUE, FALSE, EXP_REPORT);
end MODEL;
